module empty #(parameter width = 15)(
    input   [width-1 : 0] IN,
    output  [width-1 : 0] OUT
);

    // Zero Logic Module

endmodule
