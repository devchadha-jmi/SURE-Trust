module empty #(parameter width = 15)(
    input   [width-1 : 0] IN,
    input   [width-1 : 0] IN_T,
    output  [width-1 : 0] OUT,
    output  [width-1 : 0] OUT_T
);

    // Zero Logic Module

endmodule
